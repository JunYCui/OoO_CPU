`include "../define/interface.sv"

module cRAT();
/*    
input clock,
    input reset,

    sRAT_if.wr_ch wr_ch0,
    sRAT_if.wr_ch wr_ch1,   
    sRAT_if.wr_ch wr_ch2,
    sRAT_if.wr_ch wr_ch3,   

    sRAT_if.re_ch re_ch0,
    sRAT_if.re_ch re_ch1,   
    sRAT_if.re_ch re_ch2,
    sRAT_if.re_ch re_ch3, 
    sRAT_if.re_ch re_ch4,
    sRAT_if.re_ch re_ch5, 
    sRAT_if.re_ch re_ch6,
    sRAT_if.re_ch re_ch7, 

);
    
logic [8:0]cam[2**5-1:0];

    always @(posedge clock) begin
        
    end



*/
endmodule //RAT

